module top_module(clk , rst);

    input clk , rst;

    wire PCSrcE,RegWriteW,RegWriteE,ALUSrcE,MemWriteE,BranchE,RegWriteM,MemWriteM;
    wire [1:0] ResultSrcE,ResultSrcM,ResultSrcW;
    wire [2:0] ALUControlE;
    wire [4:0] RDW,RD_M,RD_W;
    wire [31:0] PCTargetE,InstrD,PCD,PCPlus4D,ResultW,RD1_E,RD2_E,Imm_Ext_E,RD_E,PCE,PCPlus4E,PCPlus4M,WriteDataM,ALU_ResultM,PCPlus4W,ALU_ResultW,ReadDataW;


    

    fetch_cycle u_fetch_cycle (
        .clk          (clk),
        .rst          (rst),
        .PCSrcE       (PCSrcE),
        .PCTargetE    (PCTargetE),
        .InstrD       (InstrD),
        .PCD          (PCD),
        .PCPlus4D     (PCPlus4D)
    );
    
    decode_cycle u_decode_cycle (
        .clk            (clk),
        .rst            (rst),
        .InstrD         (InstrD),
        .PCD            (PCD),
        .PCPlus4D       (PCPlus4D),
        .RegWriteW      (RegWriteW),
        .RDW            (RDW),
        .ResultW        (ResultW),
        .RegWriteE      (RegWriteE),
        .ALUSrcE        (ALUSrcE),
        .MemWriteE      (MemWriteE), 
        .ResultSrcE     (ResultSrcE),
        .BranchE        (BranchE),
        .ALUControlE    (ALUControlE),
        .RD1_E          (RD1_E),
        .RD2_E          (RD2_E),
        .Imm_Ext_E      (Imm_Ext_E),
        .RD_E           (RD_E),
        .PCE            (PCE),
        .PCPlus4E       (PCPlus4E),
        .RS1_E          (),
        .RS2_E          ()
    );

    execute_cycle u_execute_cycle (
        .clk            (clk),
        .rst            (rst),
        .RegWriteE      (RegWriteE),
        .ALUSrcE        (ALUSrcE),
        .MemWriteE      (MemWriteE),
        .ResultSrcE     (ResultSrcE),
        .BranchE        (BranchE),
        .ALUControlE    (ALUControlE),
        .RD1_E          (RD1_E),
        .RD2_E          (RD2_E),
        .Imm_Ext_E      (Imm_Ext_E),
        .RD_E           (RD_E),
        .PCE            (PCE),
        .PCPlus4E       (PCPlus4E),
        .PCSrcE         (PCSrcE),
        .PCTargetE      (PCTargetE),
        .RegWriteM      (RegWriteM),
        .MemWriteM      (MemWriteM),
        .ResultSrcM     (ResultSrcM),
        .RD_M           (RD_M),
        .PCPlus4M       (PCPlus4M),
        .WriteDataM     (WriteDataM),
        .ALU_ResultM    (ALU_ResultM)
    );

    memory_cycle u_memory_cycle (
        .clk            (clk),
        .rst            (rst),
        .RegWriteM      (RegWriteM),
        .MemWriteM      (MemWriteM),
        .ResultSrcM     (ResultSrcM),
        .RD_M           (RD_M),
        .PCPlus4M       (PCPlus4M),
        .WriteDataM     (WriteDataM),
        .ALU_ResultM    (ALU_ResultM),
        .RegWriteW      (RegWriteW),
        .ResultSrcW     (ResultSrcW),
        .RD_W           (RD_W),
        .PCPlus4W       (PCPlus4W),
        .ALU_ResultW    (ALU_ResultW),
        .ReadDataW      (ReadDataW)
    );

    writeback_cycle u_writeback_cycle (
        .clk            (clk),
        .rst            (rst),
        .ResultSrcW     (ResultSrcW),
        .PCPlus4W       (PCPlus4W),
        .ALU_ResultW    (ALU_ResultW),
        .ReadDataW      (ReadDataW),
        .ResultW        (ResultW)
    );




endmodule